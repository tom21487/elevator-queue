module decoder (
    input [1:0] in2,
    output [3:0] out4
);
    assign out4 = 0;
endmodule
